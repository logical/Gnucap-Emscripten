difpair ckt - simple differential pair
* modified from Spice-3 examples

*>.opt rstray cstray outwidth=80
.option method=gear

vin 1 0 sin(0 0.1 5meg) ac 1 dc 0
vcc 8 0 12
vee 9 0 -12
q1 4 2 6 0 qnl
q2 5 3 6 0 qnl
rs1 1 2 1k
rs2 3 0 1k
rc1 4 8 10k
rc2 5 8 10k
q3 6 7 9 0 qnl
q4 7 7 9 0 qnl
rbias 7 8 20k
.model qnl npn(bf=80 rb=100 va=50 tr=.4)

*>.print op v(?)
*>.op
*>.print tran qbc(q*)
*>.tran 20ns 200ns
*>.print tran cmu(q*)
*>.tran 20ns 200ns
*>.print tran vbc(q*)
*>.tran 20ns 200ns
.plot tran v(5)
*>.plot tran v(5)(2,10)
.tran 10ns 500ns

.plot ac vm(5) vp(5)
*>.plot ac vm(5)(0,100) vp(5)(-180,180)
*>.ac dec 4 10k 10ghz
.op
.ac dec 4 10k 10ghz
*>.status notime
.end
