Mesfet level 1 subthreshold characteristics
* from ngspice, modified
.param area=1.4

Vds 1 0 dc 0.1
vids 1 2 dc 0
vref 1 4 dc 0
Vgs 3 0 dc 0

z1 2 3 0 mesmod area=area
z2 4 3 0 mesmod area=1.4

.model mesmod nmf level=1 rd=46 rs=46 vt0=-1.3
+ lambda=0.03 alpha=3 beta=1.4e-3

.param area=3.5
*.print DC vids#branch
*>.print DC i(vids) i(vref)
.dc vgs -3 0 0.5

.param area=2.0
.dc vgs -3 0 0.5

.param area=1.4
.dc

.end
