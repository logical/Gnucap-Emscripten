difpair ckt - simple differential pair
* modified from Spice-3 examples

*>.opt rstray cstray phase=radians outwidth=80
.option method=gear

vin 1 0 sin(0 0.1 5meg) ac 1 dc 0
eprobe 10 0 1 0 33
vcc 8 0 12
vee 9 0 -12
q1 4 2 6 0 qnl
q2 5 3 6 0 qnl
rs1 1 2 1k
rs2 3 0 1k
rc1 4 8 10k
rc2 5 8 10k
q3 6 7 9 0 qnl
q4 7 7 9 0 qnl
rbias 7 8 20k
.model qnl npn(bf=80 rb=100 va=50 tf=4ns ptf=0)

.plot dc v(4)(-4,12) v(5)(-4,12)
.dc vin -0.2 0.2 0.01

.plot tran v(10) v(5)
*>.print tran qbe(q*)
*>.tran 10ns 300ns
*>.print tran cpi(q*)
*>.tran 10ns 300ns
*>.print tran vbe(q*)
*>.tran 10ns 300ns
*>.plot tran v(5)(2,10)
.tran 10ns 300ns

*>.print op cpi(q*)
.op

.print ac vm(5) vp(5)
*>.ac dec 5 10k 1ghz
.plot ac vm(5)
.plot ac vp(5)
*>.plot ac vm(5)(0,100) vp(5)(-2,2)
.ac dec 5 10k 1ghz
.status notime
.end
